module D_FF(D, clk, rst, q);  wire _0_;  input D;  input clk;  output q;  input rst;  AND2X2 _1_ (    .A(D),    .B(rst),    .Y(_0_)  );  DFFPOSX1 _2_ (    .CLK(clk),    .D(_0_),    .Q(q)  );endmodulemodule simpleR_R(a, d, clk, rst, y);  input a;  wire c;  input clk;  input d;  wire g;  input rst;  output y;  OR2X2 _0_ (    .A(c),    .B(a),    .Y(g)  );  D_FF dff1 (    .D(d),    .clk(clk),    .q(c),    .rst(rst)  );  D_FF dff2 (    .D(g),    .clk(clk),    .q(y),    .rst(rst)  );endmodule
