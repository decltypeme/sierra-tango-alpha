// // file: test.v
// // author: @hussama

// `timescale 1ns/1ns

// module mux4_1(
    // output [3:0] out,
    // input [3:0] x,
    // input [3:0] y,
    // input  sel
    // );

// assign out= (sel==1'b0)? x:
				     // y;
// endmodule

// module fourbitmux2X1ToRegToReg(output [3:0] out,
    // input [3:0] x,
    // input [3:0] y,
    // input  sel,
    // input clk);
    
    // wire [3:0] imm;
    
    // mux4_1 _mux4_1(imm,x,y,sel);
    
    // reg [3:0] r1;
    // reg [3:0] r2;
        
    // always @(posedge clk)
    // begin
        // r1 <= imm;
        // r2 <= r1;
    // end
    
    // assign out = r2; 

// endmodule

/* Generated by Yosys 0.6 (git sha1 UNKNOWN, clang 3.4-1ubuntu3 -fPIC -Os) */

module fourbitmux2X1ToRegToReg(out, x, y, sel, clk);
  input clk;
  wire [3:0] imm;
  output [3:0] out;
  wire [3:0] r1;
  input sel;
  input [3:0] x;
  input [3:0] y;
  DFFPOSX1 _0_ (
    .CLK(clk),
    .D(r1[0]),
    .Q(out[0])
  );
  DFFPOSX1 _1_ (
    .CLK(clk),
    .D(r1[1]),
    .Q(out[1])
  );
  DFFPOSX1 _2_ (
    .CLK(clk),
    .D(r1[2]),
    .Q(out[2])
  );
  DFFPOSX1 _3_ (
    .CLK(clk),
    .D(r1[3]),
    .Q(out[3])
  );
  DFFPOSX1 _4_ (
    .CLK(clk),
    .D(imm[0]),
    .Q(r1[0])
  );
  DFFPOSX1 _5_ (
    .CLK(clk),
    .D(imm[1]),
    .Q(r1[1])
  );
  DFFPOSX1 _6_ (
    .CLK(clk),
    .D(imm[2]),
    .Q(r1[2])
  );
  DFFPOSX1 _7_ (
    .CLK(clk),
    .D(imm[3]),
    .Q(r1[3])
  );
  mux4_1 _mux4_1 (
    .out(imm),
    .sel(sel),
    .x(x),
    .y(y)
  );
endmodule

module mux4_1(out, x, y, sel);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  output [3:0] out;
  input sel;
  input [3:0] x;
  input [3:0] y;
  INVX1 _08_ (
    .A(x[0]),
    .Y(_00_)
  );
  NAND2X1 _09_ (
    .A(y[0]),
    .B(sel),
    .Y(_01_)
  );
  OAI21X1 _10_ (
    .A(sel),
    .B(_00_),
    .C(_01_),
    .Y(out[0])
  );
  INVX1 _11_ (
    .A(x[1]),
    .Y(_02_)
  );
  NAND2X1 _12_ (
    .A(sel),
    .B(y[1]),
    .Y(_03_)
  );
  OAI21X1 _13_ (
    .A(sel),
    .B(_02_),
    .C(_03_),
    .Y(out[1])
  );
  INVX1 _14_ (
    .A(x[2]),
    .Y(_04_)
  );
  NAND2X1 _15_ (
    .A(sel),
    .B(y[2]),
    .Y(_05_)
  );
  OAI21X1 _16_ (
    .A(sel),
    .B(_04_),
    .C(_05_),
    .Y(out[2])
  );
  INVX1 _17_ (
    .A(x[3]),
    .Y(_06_)
  );
  NAND2X1 _18_ (
    .A(sel),
    .B(y[3]),
    .Y(_07_)
  );
  OAI21X1 _19_ (
    .A(sel),
    .B(_06_),
    .C(_07_),
    .Y(out[3])
  );
endmodule

