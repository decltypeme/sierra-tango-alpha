module bits(a, b); input a; output b; INVX1 _0_ ( .A(a), .Y(b) );endmodule
